
module delta (    
    input reg [4:0] data,
    input reg [4:0] threshold,
    input reg [4:0] prev,
    input wire off_spike,
    output wire spike[1:0]
);

// compares the difference between current data and previous against a threshold

endmodule

